module rnn_recurrent();

	logic [15:0] R[0:31][0:31];

	assign R[0][0]  = 16'b0000000001001111;
	assign R[0][1]  = 16'b0000000001110001;
	assign R[0][2]  = 16'b1111111110010000;
	assign R[0][3]  = 16'b0000000000101000;
	assign R[0][4]  = 16'b0000000001000010;
	assign R[0][5]  = 16'b1111111111011110;
	assign R[0][6]  = 16'b0000000001101001;
	assign R[0][7]  = 16'b0000000010110000;
	assign R[0][8]  = 16'b0000000001001110;
	assign R[0][9]  = 16'b1111111111110110;
	assign R[0][10] = 16'b1111111110110101;
	assign R[0][11] = 16'b1111111111000010;
	assign R[0][12] = 16'b0000000001001100;
	assign R[0][13] = 16'b0000000000100011;
	assign R[0][14] = 16'b0000000000001100;
	assign R[0][15] = 16'b0000000100110001;
	assign R[0][16] = 16'b1111111111010100;
	assign R[0][17] = 16'b0000000000001101;
	assign R[0][18] = 16'b1111111111101100;
	assign R[0][19] = 16'b0000000000000011;
	assign R[0][20] = 16'b0000000000011100;
	assign R[0][21] = 16'b1111111111110101;
	assign R[0][22] = 16'b0000000000011011;
	assign R[0][23] = 16'b1111111111101110;
	assign R[0][24] = 16'b1111111110110011;
	assign R[0][25] = 16'b0000000000010010;
	assign R[0][26] = 16'b1111111111000000;
	assign R[0][27] = 16'b1111111111001110;
	assign R[0][28] = 16'b1111111101100111;
	assign R[0][29] = 16'b0000000000001011;
	assign R[0][30] = 16'b0000000000000010;
	assign R[0][31] = 16'b1111111111011101;
	assign R[1][0]  = 16'b0000000000100010;
	assign R[1][1]  = 16'b0000000001111101;
	assign R[1][2]  = 16'b0000000000011101;
	assign R[1][3]  = 16'b1111111111010011;
	assign R[1][4]  = 16'b0000000001010000;
	assign R[1][5]  = 16'b1111111111100000;
	assign R[1][6]  = 16'b0000000000000100;
	assign R[1][7]  = 16'b1111111110101010;
	assign R[1][8]  = 16'b0000000000101111;
	assign R[1][9]  = 16'b0000000001011000;
	assign R[1][10] = 16'b1111111111110011;
	assign R[1][11] = 16'b1111111111011011;
	assign R[1][12] = 16'b0000000001010100;
	assign R[1][13] = 16'b0000000000101100;
	assign R[1][14] = 16'b1111111110010111;
	assign R[1][15] = 16'b0000000000101111;
	assign R[1][16] = 16'b1111111110011010;
	assign R[1][17] = 16'b0000000001110000;
	assign R[1][18] = 16'b1111111101100111;
	assign R[1][19] = 16'b1111111111110000;
	assign R[1][20] = 16'b1111111111101001;
	assign R[1][21] = 16'b1111111111011110;
	assign R[1][22] = 16'b1111111111101110;
	assign R[1][23] = 16'b0000000000001101;
	assign R[1][24] = 16'b0000000000010001;
	assign R[1][25] = 16'b1111111111101110;
	assign R[1][26] = 16'b1111111110110100;
	assign R[1][27] = 16'b1111111111101101;
	assign R[1][28] = 16'b0000000001000101;
	assign R[1][29] = 16'b1111111111110001;
	assign R[1][30] = 16'b0000000000010101;
	assign R[1][31] = 16'b0000000000011000;
	assign R[2][0]  = 16'b1111111111101011;
	assign R[2][1]  = 16'b0000000010111001;
	assign R[2][2]  = 16'b0000000000100110;
	assign R[2][3]  = 16'b1111111111101110;
	assign R[2][4]  = 16'b0000000000000000;
	assign R[2][5]  = 16'b1111111111100001;
	assign R[2][6]  = 16'b1111111111011000;
	assign R[2][7]  = 16'b1111111110101010;
	assign R[2][8]  = 16'b0000000000011010;
	assign R[2][9]  = 16'b1111111110111001;
	assign R[2][10] = 16'b0000000001001111;
	assign R[2][11] = 16'b0000000000010111;
	assign R[2][12] = 16'b1111111110110001;
	assign R[2][13] = 16'b0000000000000000;
	assign R[2][14] = 16'b0000000000110011;
	assign R[2][15] = 16'b0000000010010110;
	assign R[2][16] = 16'b0000000000001011;
	assign R[2][17] = 16'b0000000010001000;
	assign R[2][18] = 16'b0000000000000000;
	assign R[2][19] = 16'b0000000000010111;
	assign R[2][20] = 16'b1111111111011010;
	assign R[2][21] = 16'b1111111101110110;
	assign R[2][22] = 16'b0000000000010110;
	assign R[2][23] = 16'b0000000001111100;
	assign R[2][24] = 16'b1111111111111100;
	assign R[2][25] = 16'b0000000000000001;
	assign R[2][26] = 16'b1111111111101001;
	assign R[2][27] = 16'b0000000000000010;
	assign R[2][28] = 16'b0000000001001001;
	assign R[2][29] = 16'b0000000001100110;
	assign R[2][30] = 16'b0000000000000111;
	assign R[2][31] = 16'b0000000101001011;
	assign R[3][0]  = 16'b0000000000000110;
	assign R[3][1]  = 16'b0000000000000000;
	assign R[3][2]  = 16'b0000000000101001;
	assign R[3][3]  = 16'b0000000010000011;
	assign R[3][4]  = 16'b0000000000001011;
	assign R[3][5]  = 16'b1111111110111111;
	assign R[3][6]  = 16'b0000000001001110;
	assign R[3][7]  = 16'b0000000000001110;
	assign R[3][8]  = 16'b0000000000010111;
	assign R[3][9]  = 16'b0000000000110111;
	assign R[3][10] = 16'b1111111111100000;
	assign R[3][11] = 16'b1111111111011100;
	assign R[3][12] = 16'b0000000001001111;
	assign R[3][13] = 16'b0000000000110000;
	assign R[3][14] = 16'b1111111111111100;
	assign R[3][15] = 16'b1111111111101100;
	assign R[3][16] = 16'b0000000000000110;
	assign R[3][17] = 16'b1111111110100001;
	assign R[3][18] = 16'b0000000000010101;
	assign R[3][19] = 16'b1111111110101111;
	assign R[3][20] = 16'b1111111111111001;
	assign R[3][21] = 16'b1111111111111001;
	assign R[3][22] = 16'b1111111111110010;
	assign R[3][23] = 16'b1111111111001100;
	assign R[3][24] = 16'b0000000001110101;
	assign R[3][25] = 16'b1111111111111110;
	assign R[3][26] = 16'b1111111111100100;
	assign R[3][27] = 16'b0000000000010110;
	assign R[3][28] = 16'b1111111110101100;
	assign R[3][29] = 16'b0000000001011110;
	assign R[3][30] = 16'b0000000000000100;
	assign R[3][31] = 16'b1111111110100011;
	assign R[4][0]  = 16'b0000000000001101;
	assign R[4][1]  = 16'b0000000001101111;
	assign R[4][2]  = 16'b0000000000000011;
	assign R[4][3]  = 16'b1111111111100000;
	assign R[4][4]  = 16'b1111111110101001;
	assign R[4][5]  = 16'b1111111111101010;
	assign R[4][6]  = 16'b1111111110000100;
	assign R[4][7]  = 16'b1111111110101001;
	assign R[4][8]  = 16'b1111111110101000;
	assign R[4][9]  = 16'b1111111110010010;
	assign R[4][10] = 16'b0000000000010000;
	assign R[4][11] = 16'b1111111111101010;
	assign R[4][12] = 16'b0000000011001101;
	assign R[4][13] = 16'b0000000000100010;
	assign R[4][14] = 16'b0000000000110110;
	assign R[4][15] = 16'b1111111101000110;
	assign R[4][16] = 16'b0000000000110110;
	assign R[4][17] = 16'b0000000000001110;
	assign R[4][18] = 16'b0000000000001011;
	assign R[4][19] = 16'b0000000000100000;
	assign R[4][20] = 16'b0000000000001010;
	assign R[4][21] = 16'b1111111111111100;
	assign R[4][22] = 16'b0000000000111100;
	assign R[4][23] = 16'b0000000000111000;
	assign R[4][24] = 16'b1111111110101011;
	assign R[4][25] = 16'b0000000000111100;
	assign R[4][26] = 16'b0000000000111000;
	assign R[4][27] = 16'b1111111110011010;
	assign R[4][28] = 16'b1111111111001010;
	assign R[4][29] = 16'b0000000001000101;
	assign R[4][30] = 16'b0000000000010111;
	assign R[4][31] = 16'b1111111111101000;
	assign R[5][0]  = 16'b0000000000010100;
	assign R[5][1]  = 16'b1111111110100000;
	assign R[5][2]  = 16'b1111111101111000;
	assign R[5][3]  = 16'b1111111111010101;
	assign R[5][4]  = 16'b0000000001100011;
	assign R[5][5]  = 16'b0000000010000100;
	assign R[5][6]  = 16'b0000000001100111;
	assign R[5][7]  = 16'b0000000001101001;
	assign R[5][8]  = 16'b0000000001010001;
	assign R[5][9]  = 16'b1111111111100000;
	assign R[5][10] = 16'b0000000001100100;
	assign R[5][11] = 16'b1111111110000111;
	assign R[5][12] = 16'b1111111110010101;
	assign R[5][13] = 16'b0000000000111001;
	assign R[5][14] = 16'b1111111111010101;
	assign R[5][15] = 16'b0000000001011010;
	assign R[5][16] = 16'b0000000000001100;
	assign R[5][17] = 16'b1111111100101111;
	assign R[5][18] = 16'b1111111110101100;
	assign R[5][19] = 16'b1111111111110001;
	assign R[5][20] = 16'b0000000000010100;
	assign R[5][21] = 16'b0000000000111001;
	assign R[5][22] = 16'b0000000001001110;
	assign R[5][23] = 16'b0000000001001100;
	assign R[5][24] = 16'b1111111110001101;
	assign R[5][25] = 16'b0000000000111010;
	assign R[5][26] = 16'b1111111111000000;
	assign R[5][27] = 16'b1111111110100101;
	assign R[5][28] = 16'b0000000000001111;
	assign R[5][29] = 16'b0000000001010111;
	assign R[5][30] = 16'b1111111111000101;
	assign R[5][31] = 16'b0000000100001100;
	assign R[6][0]  = 16'b0000000001100100;
	assign R[6][1]  = 16'b1111111110101000;
	assign R[6][2]  = 16'b0000000000000001;
	assign R[6][3]  = 16'b1111111110011111;
	assign R[6][4]  = 16'b0000000001011011;
	assign R[6][5]  = 16'b0000000000000100;
	assign R[6][6]  = 16'b0000000000101010;
	assign R[6][7]  = 16'b0000000001001101;
	assign R[6][8]  = 16'b0000000001000001;
	assign R[6][9]  = 16'b0000000000011101;
	assign R[6][10] = 16'b0000000000100101;
	assign R[6][11] = 16'b1111111111001010;
	assign R[6][12] = 16'b0000000000010001;
	assign R[6][13] = 16'b0000000000101100;
	assign R[6][14] = 16'b1111111111010110;
	assign R[6][15] = 16'b0000000001001001;
	assign R[6][16] = 16'b1111111110111011;
	assign R[6][17] = 16'b1111111111010010;
	assign R[6][18] = 16'b1111111101110100;
	assign R[6][19] = 16'b0000000001110101;
	assign R[6][20] = 16'b1111111111110111;
	assign R[6][21] = 16'b0000000000110110;
	assign R[6][22] = 16'b0000000001000011;
	assign R[6][23] = 16'b0000000000111011;
	assign R[6][24] = 16'b1111111110111111;
	assign R[6][25] = 16'b1111111111010111;
	assign R[6][26] = 16'b0000000000010011;
	assign R[6][27] = 16'b0000000000010111;
	assign R[6][28] = 16'b1111111111100000;
	assign R[6][29] = 16'b0000000001001100;
	assign R[6][30] = 16'b0000000000000100;
	assign R[6][31] = 16'b0000000001000111;
	assign R[7][0]  = 16'b0000000000000000;
	assign R[7][1]  = 16'b0000000000001000;
	assign R[7][2]  = 16'b0000000011001101;
	assign R[7][3]  = 16'b1111111111000110;
	assign R[7][4]  = 16'b1111111111101110;
	assign R[7][5]  = 16'b0000000000001110;
	assign R[7][6]  = 16'b0000000010000110;
	assign R[7][7]  = 16'b0000000000110111;
	assign R[7][8]  = 16'b1111111111001111;
	assign R[7][9]  = 16'b1111111111011011;
	assign R[7][10] = 16'b0000000000001100;
	assign R[7][11] = 16'b0000000001100011;
	assign R[7][12] = 16'b1111111111010101;
	assign R[7][13] = 16'b0000000000000111;
	assign R[7][14] = 16'b0000000001010110;
	assign R[7][15] = 16'b0000000110011100;
	assign R[7][16] = 16'b1111111111100100;
	assign R[7][17] = 16'b1111111110111110;
	assign R[7][18] = 16'b0000000001000100;
	assign R[7][19] = 16'b0000000000011100;
	assign R[7][20] = 16'b0000000000001000;
	assign R[7][21] = 16'b1111111111101111;
	assign R[7][22] = 16'b0000000000011011;
	assign R[7][23] = 16'b1111111101110101;
	assign R[7][24] = 16'b0000000000111011;
	assign R[7][25] = 16'b1111111111101001;
	assign R[7][26] = 16'b0000000000001110;
	assign R[7][27] = 16'b1111111111010101;
	assign R[7][28] = 16'b0000000001101001;
	assign R[7][29] = 16'b0000000000110110;
	assign R[7][30] = 16'b0000000001010001;
	assign R[7][31] = 16'b0000000000110010;
	assign R[8][0]  = 16'b0000000010010110;
	assign R[8][1]  = 16'b0000000000111111;
	assign R[8][2]  = 16'b1111111111001011;
	assign R[8][3]  = 16'b1111111111111010;
	assign R[8][4]  = 16'b0000000000011110;
	assign R[8][5]  = 16'b0000000001101010;
	assign R[8][6]  = 16'b1111111110001111;
	assign R[8][7]  = 16'b0000000001011100;
	assign R[8][8]  = 16'b0000000000011111;
	assign R[8][9]  = 16'b0000000001010101;
	assign R[8][10] = 16'b0000000001001110;
	assign R[8][11] = 16'b1111111111010110;
	assign R[8][12] = 16'b1111111110001101;
	assign R[8][13] = 16'b1111111110110000;
	assign R[8][14] = 16'b1111111111101110;
	assign R[8][15] = 16'b0000000001110100;
	assign R[8][16] = 16'b1111111111001000;
	assign R[8][17] = 16'b1111111111010000;
	assign R[8][18] = 16'b1111111101010100;
	assign R[8][19] = 16'b1111111110110111;
	assign R[8][20] = 16'b0000000000010001;
	assign R[8][21] = 16'b1111111110100100;
	assign R[8][22] = 16'b0000000000001000;
	assign R[8][23] = 16'b0000000000001010;
	assign R[8][24] = 16'b0000000010000101;
	assign R[8][25] = 16'b0000000000011000;
	assign R[8][26] = 16'b0000000001000111;
	assign R[8][27] = 16'b0000000010100010;
	assign R[8][28] = 16'b1111111111000100;
	assign R[8][29] = 16'b1111111110111011;
	assign R[8][30] = 16'b1111111110111000;
	assign R[8][31] = 16'b0000000001000001;
	assign R[9][0]  = 16'b0000000000010011;
	assign R[9][1]  = 16'b1111111110111001;
	assign R[9][2]  = 16'b1111111111110111;
	assign R[9][3]  = 16'b1111111111001100;
	assign R[9][4]  = 16'b0000000000110000;
	assign R[9][5]  = 16'b1111111110011101;
	assign R[9][6]  = 16'b1111111110110001;
	assign R[9][7]  = 16'b1111111111000011;
	assign R[9][8]  = 16'b1111111110110111;
	assign R[9][9]  = 16'b0000000011000110;
	assign R[9][10] = 16'b1111111111001101;
	assign R[9][11] = 16'b1111111110111101;
	assign R[9][12] = 16'b1111111101001011;
	assign R[9][13] = 16'b0000000000010101;
	assign R[9][14] = 16'b1111111111011111;
	assign R[9][15] = 16'b1111111101011101;
	assign R[9][16] = 16'b1111111111100001;
	assign R[9][17] = 16'b0000000000011001;
	assign R[9][18] = 16'b1111111110111111;
	assign R[9][19] = 16'b0000000000000000;
	assign R[9][20] = 16'b0000000000001100;
	assign R[9][21] = 16'b0000000000000000;
	assign R[9][22] = 16'b0000000000010111;
	assign R[9][23] = 16'b1111111111110111;
	assign R[9][24] = 16'b0000000001001010;
	assign R[9][25] = 16'b1111111111110111;
	assign R[9][26] = 16'b1111111110011001;
	assign R[9][27] = 16'b0000000001000100;
	assign R[9][28] = 16'b0000000000110110;
	assign R[9][29] = 16'b0000000010001011;
	assign R[9][30] = 16'b1111111110111010;
	assign R[9][31] = 16'b1111111101111100;
	assign R[10][0] = 16'b0000000000011101;
	assign R[10][1] = 16'b1111111110010011;
	assign R[10][2] = 16'b0000000000001111;
	assign R[10][3] = 16'b1111111110000001;
	assign R[10][4] = 16'b1111111111001111;
	assign R[10][5] = 16'b0000000000100010;
	assign R[10][6] = 16'b1111111111100010;
	assign R[10][7] = 16'b0000000000100010;
	assign R[10][8] = 16'b0000000001010001;
	assign R[10][9] = 16'b0000000010011011;
	assign R[10][10] = 16'b1111111110110100;
	assign R[10][11] = 16'b1111111111011000;
	assign R[10][12] = 16'b0000000010010011;
	assign R[10][13] = 16'b0000000000100100;
	assign R[10][14] = 16'b1111111111111100;
	assign R[10][15] = 16'b1111111111111110;
	assign R[10][16] = 16'b0000000000111001;
	assign R[10][17] = 16'b0000000010101111;
	assign R[10][18] = 16'b1111111101111111;
	assign R[10][19] = 16'b0000000000100100;
	assign R[10][20] = 16'b0000000000111011;
	assign R[10][21] = 16'b0000000001010010;
	assign R[10][22] = 16'b0000000001101001;
	assign R[10][23] = 16'b0000000000011100;
	assign R[10][24] = 16'b0000000000100100;
	assign R[10][25] = 16'b1111111101001010;
	assign R[10][26] = 16'b1111111110101011;
	assign R[10][27] = 16'b0000000001101101;
	assign R[10][28] = 16'b1111111110110111;
	assign R[10][29] = 16'b1111111111111100;
	assign R[10][30] = 16'b0000000000001101;
	assign R[10][31] = 16'b0000000000001001;
	assign R[11][0]  = 16'b1111111101010010;
	assign R[11][1]  = 16'b0000000000010001;
	assign R[11][2]  = 16'b0000000000000110;
	assign R[11][3]  = 16'b0000000000110000;
	assign R[11][4]  = 16'b0000000000100110;
	assign R[11][5]  = 16'b0000000001011000;
	assign R[11][6]  = 16'b1111111101111001;
	assign R[11][7]  = 16'b0000000010010100;
	assign R[11][8]  = 16'b0000000000111010;
	assign R[11][9]  = 16'b0000000000001101;
	assign R[11][10] = 16'b0000000001000000;
	assign R[11][11] = 16'b0000000001000111;
	assign R[11][12] = 16'b0000000001111000;
	assign R[11][13] = 16'b1111111111100001;
	assign R[11][14] = 16'b1111111111001111;
	assign R[11][15] = 16'b1111111110111110;
	assign R[11][16] = 16'b0000000001000101;
	assign R[11][17] = 16'b0000000001100011;
	assign R[11][18] = 16'b0000000000101011;
	assign R[11][19] = 16'b1111111110011011;
	assign R[11][20] = 16'b0000000000111001;
	assign R[11][21] = 16'b0000000000001111;
	assign R[11][22] = 16'b0000000000100101;
	assign R[11][23] = 16'b0000000001011001;
	assign R[11][24] = 16'b0000000000100001;
	assign R[11][25] = 16'b0000000000100101;
	assign R[11][26] = 16'b1111111111101010;
	assign R[11][27] = 16'b1111111011101111;
	assign R[11][28] = 16'b1111111111111010;
	assign R[11][29] = 16'b1111111111001010;
	assign R[11][30] = 16'b1111111111101110;
	assign R[11][31] = 16'b0000000001000000;
	assign R[12][0]  = 16'b1111111111011110;
	assign R[12][1]  = 16'b1111111111110000;
	assign R[12][2]  = 16'b1111111111011010;
	assign R[12][3]  = 16'b0000000000100110;
	assign R[12][4]  = 16'b1111111111000001;
	assign R[12][5]  = 16'b0000000000011111;
	assign R[12][6]  = 16'b0000000000101100;
	assign R[12][7]  = 16'b1111111100111110;
	assign R[12][8]  = 16'b1111111111011010;
	assign R[12][9]  = 16'b1111111111001101;
	assign R[12][10] = 16'b0000000000001010;
	assign R[12][11] = 16'b0000000000101010;
	assign R[12][12] = 16'b0000000001100001;
	assign R[12][13] = 16'b1111111111101000;
	assign R[12][14] = 16'b1111111111100100;
	assign R[12][15] = 16'b0000000100111110;
	assign R[12][16] = 16'b1111111110111111;
	assign R[12][17] = 16'b1111111101110000;
	assign R[12][18] = 16'b1111111111000100;
	assign R[12][19] = 16'b0000000000100011;
	assign R[12][20] = 16'b0000000000110011;
	assign R[12][21] = 16'b1111111111100011;
	assign R[12][22] = 16'b0000000010000101;
	assign R[12][23] = 16'b1111111111101001;
	assign R[12][24] = 16'b1111111111010111;
	assign R[12][25] = 16'b1111111111100001;
	assign R[12][26] = 16'b0000000000111000;
	assign R[12][27] = 16'b0000000001000011;
	assign R[12][28] = 16'b0000000000100111;
	assign R[12][29] = 16'b0000000000000011;
	assign R[12][30] = 16'b1111111111110101;
	assign R[12][31] = 16'b1111111110101101;
	assign R[13][0]  = 16'b1111111101111111;
	assign R[13][1]  = 16'b0000000001111010;
	assign R[13][2]  = 16'b1111111110010001;
	assign R[13][3]  = 16'b0000000000100101;
	assign R[13][4]  = 16'b0000000000010110;
	assign R[13][5]  = 16'b1111111111110101;
	assign R[13][6]  = 16'b1111111110001010;
	assign R[13][7]  = 16'b0000000000100010;
	assign R[13][8]  = 16'b1111111111101101;
	assign R[13][9]  = 16'b1111111111001110;
	assign R[13][10] = 16'b1111111111010101;
	assign R[13][11] = 16'b1111111111001010;
	assign R[13][12] = 16'b1111111110100110;
	assign R[13][13] = 16'b0000000000010010;
	assign R[13][14] = 16'b1111111111110110;
	assign R[13][15] = 16'b1111111111110001;
	assign R[13][16] = 16'b0000000000001101;
	assign R[13][17] = 16'b0000000010000111;
	assign R[13][18] = 16'b1111111101100000;
	assign R[13][19] = 16'b0000000000011010;
	assign R[13][20] = 16'b0000000000000001;
	assign R[13][21] = 16'b0000000000011001;
	assign R[13][22] = 16'b1111111110001010;
	assign R[13][23] = 16'b1111111111110010;
	assign R[13][24] = 16'b1111111111000010;
	assign R[13][25] = 16'b0000000000010011;
	assign R[13][26] = 16'b1111111111101010;
	assign R[13][27] = 16'b1111111111000000;
	assign R[13][28] = 16'b0000000000101100;
	assign R[13][29] = 16'b1111111111101111;
	assign R[13][30] = 16'b1111111111011011;
	assign R[13][31] = 16'b1111111110001110;
	assign R[14][0]  = 16'b0000000000010111;
	assign R[14][1]  = 16'b0000000000010010;
	assign R[14][2]  = 16'b1111111111100100;
	assign R[14][3]  = 16'b1111111111110010;
	assign R[14][4]  = 16'b1111111111011011;
	assign R[14][5]  = 16'b0000000001110001;
	assign R[14][6]  = 16'b0000000001001100;
	assign R[14][7]  = 16'b0000000010011010;
	assign R[14][8]  = 16'b0000000001111111;
	assign R[14][9]  = 16'b1111111111111010;
	assign R[14][10] = 16'b1111111110000100;
	assign R[14][11] = 16'b0000000000010001;
	assign R[14][12] = 16'b0000000000101000;
	assign R[14][13] = 16'b0000000001010011;
	assign R[14][14] = 16'b0000000100101000;
	assign R[14][15] = 16'b1111111101101100;
	assign R[14][16] = 16'b1111111110100101;
	assign R[14][17] = 16'b0000000001111000;
	assign R[14][18] = 16'b0000000001000111;
	assign R[14][19] = 16'b0000000000100011;
	assign R[14][20] = 16'b0000000001101100;
	assign R[14][21] = 16'b0000000001000001;
	assign R[14][22] = 16'b0000000001000001;
	assign R[14][23] = 16'b1111111111101100;
	assign R[14][24] = 16'b1111111110001110;
	assign R[14][25] = 16'b0000000000111110;
	assign R[14][26] = 16'b1111111101101110;
	assign R[14][27] = 16'b1111111101100011;
	assign R[14][28] = 16'b0000000000011100;
	assign R[14][29] = 16'b0000000001110111;
	assign R[14][30] = 16'b1111111110001011;
	assign R[14][31] = 16'b0000000001101101;
	assign R[15][0]  = 16'b1111111111111111;
	assign R[15][1]  = 16'b0000000000110001;
	assign R[15][2]  = 16'b1111111101101100;
	assign R[15][3]  = 16'b1111111110000110;
	assign R[15][4]  = 16'b0000000000001001;
	assign R[15][5]  = 16'b0000000001000001;
	assign R[15][6]  = 16'b0000000001100111;
	assign R[15][7]  = 16'b1111111111111101;
	assign R[15][8]  = 16'b0000000000010101;
	assign R[15][9]  = 16'b0000000000110000;
	assign R[15][10] = 16'b1111111110010101;
	assign R[15][11] = 16'b1111111111100110;
	assign R[15][12] = 16'b1111111110101101;
	assign R[15][13] = 16'b0000000001001010;
	assign R[15][14] = 16'b1111111111011101;
	assign R[15][15] = 16'b0000000100001100;
	assign R[15][16] = 16'b1111111101010111;
	assign R[15][17] = 16'b0000000001000101;
	assign R[15][18] = 16'b0000000000010110;
	assign R[15][19] = 16'b0000000001001000;
	assign R[15][20] = 16'b0000000000011100;
	assign R[15][21] = 16'b0000000000001110;
	assign R[15][22] = 16'b0000000000010000;
	assign R[15][23] = 16'b0000000001100011;
	assign R[15][24] = 16'b1111111111100000;
	assign R[15][25] = 16'b1111111100111000;
	assign R[15][26] = 16'b0000000000001001;
	assign R[15][27] = 16'b1111111110000100;
	assign R[15][28] = 16'b1111111111011110;
	assign R[15][29] = 16'b0000000001000011;
	assign R[15][30] = 16'b1111111111000000;
	assign R[15][31] = 16'b0000000010100110;
	assign R[16][0]  = 16'b1111111111101001;
	assign R[16][1]  = 16'b0000000000010101;
	assign R[16][2]  = 16'b1111111111011010;
	assign R[16][3]  = 16'b1111111111000001;
	assign R[16][4]  = 16'b0000000000110010;
	assign R[16][5]  = 16'b0000000000011111;
	assign R[16][6]  = 16'b1111111111110101;
	assign R[16][7]  = 16'b0000000000011000;
	assign R[16][8]  = 16'b1111111110110000;
	assign R[16][9]  = 16'b0000000001010100;
	assign R[16][10] = 16'b0000000000010001;
	assign R[16][11] = 16'b1111111110100100;
	assign R[16][12] = 16'b1111111100100110;
	assign R[16][13] = 16'b1111111111010000;
	assign R[16][14] = 16'b0000000001101000;
	assign R[16][15] = 16'b1111111110111010;
	assign R[16][16] = 16'b1111111111110110;
	assign R[16][17] = 16'b0000000000000000;
	assign R[16][18] = 16'b1111111111101000;
	assign R[16][19] = 16'b1111111111010101;
	assign R[16][20] = 16'b0000000001010111;
	assign R[16][21] = 16'b1111111110011100;
	assign R[16][22] = 16'b1111111110011011;
	assign R[16][23] = 16'b1111111110111100;
	assign R[16][24] = 16'b0000000000011001;
	assign R[16][25] = 16'b1111111111000111;
	assign R[16][26] = 16'b0000000000011001;
	assign R[16][27] = 16'b0000000000100110;
	assign R[16][28] = 16'b1111111111100110;
	assign R[16][29] = 16'b1111111111000001;
	assign R[16][30] = 16'b0000000000000000;
	assign R[16][31] = 16'b0000000001010100;
	assign R[17][0]  = 16'b0000000000000111;
	assign R[17][1]  = 16'b1111111110101000;
	assign R[17][2]  = 16'b0000000000010100;
	assign R[17][3]  = 16'b0000000000011101;
	assign R[17][4]  = 16'b1111111101111001;
	assign R[17][5]  = 16'b1111111111100001;
	assign R[17][6]  = 16'b0000000000101011;
	assign R[17][7]  = 16'b1111111111110100;
	assign R[17][8]  = 16'b1111111111011001;
	assign R[17][9]  = 16'b0000000000101001;
	assign R[17][10] = 16'b0000000000001010;
	assign R[17][11] = 16'b1111111111101101;
	assign R[17][12] = 16'b1111111111011111;
	assign R[17][13] = 16'b0000000000011000;
	assign R[17][14] = 16'b1111111111100001;
	assign R[17][15] = 16'b0000000001101101;
	assign R[17][16] = 16'b0000000000110011;
	assign R[17][17] = 16'b1111111110111010;
	assign R[17][18] = 16'b0000000001100111;
	assign R[17][19] = 16'b1111111111100100;
	assign R[17][20] = 16'b1111111111011110;
	assign R[17][21] = 16'b1111111110110110;
	assign R[17][22] = 16'b0000000001001111;
	assign R[17][23] = 16'b1111111111011010;
	assign R[17][24] = 16'b0000000001001110;
	assign R[17][25] = 16'b0000000000111111;
	assign R[17][26] = 16'b0000000000110001;
	assign R[17][27] = 16'b0000000000101011;
	assign R[17][28] = 16'b0000000000110101;
	assign R[17][29] = 16'b1111111110110001;
	assign R[17][30] = 16'b0000000001011001;
	assign R[17][31] = 16'b0000000010010101;
	assign R[18][0]  = 16'b1111111111110101;
	assign R[18][1]  = 16'b0000000000111101;
	assign R[18][2]  = 16'b1111111110110001;
	assign R[18][3]  = 16'b0000000000101001;
	assign R[18][4]  = 16'b0000000000011000;
	assign R[18][5]  = 16'b0000000001000100;
	assign R[18][6]  = 16'b1111111011100100;
	assign R[18][7]  = 16'b1111111111101011;
	assign R[18][8]  = 16'b1111111110111110;
	assign R[18][9]  = 16'b1111111111110111;
	assign R[18][10] = 16'b0000000000101011;
	assign R[18][11] = 16'b0000000000100010;
	assign R[18][12] = 16'b0000000000100001;
	assign R[18][13] = 16'b0000000000010000;
	assign R[18][14] = 16'b1111111111001100;
	assign R[18][15] = 16'b0000000010111100;
	assign R[18][16] = 16'b0000000000011111;
	assign R[18][17] = 16'b1111111111111011;
	assign R[18][18] = 16'b1111111111110011;
	assign R[18][19] = 16'b0000000011010100;
	assign R[18][20] = 16'b0000000001100000;
	assign R[18][21] = 16'b0000000000011101;
	assign R[18][22] = 16'b0000000000000011;
	assign R[18][23] = 16'b1111111111010111;
	assign R[18][24] = 16'b0000000001000001;
	assign R[18][25] = 16'b1111111111111001;
	assign R[18][26] = 16'b1111111111111110;
	assign R[18][27] = 16'b1111111111101111;
	assign R[18][28] = 16'b1111111110010101;
	assign R[18][29] = 16'b0000000000000100;
	assign R[18][30] = 16'b1111111111110110;
	assign R[18][31] = 16'b1111111100101100;
	assign R[19][0]  = 16'b1111111111101100;
	assign R[19][1]  = 16'b1111111110111010;
	assign R[19][2]  = 16'b1111111111011010;
	assign R[19][3]  = 16'b1111111110101111;
	assign R[19][4]  = 16'b0000000001001100;
	assign R[19][5]  = 16'b1111111111101101;
	assign R[19][6]  = 16'b0000000100101010;
	assign R[19][7]  = 16'b0000000000101011;
	assign R[19][8]  = 16'b0000000000001111;
	assign R[19][9]  = 16'b0000000000100001;
	assign R[19][10] = 16'b0000000000101111;
	assign R[19][11] = 16'b1111111110000010;
	assign R[19][12] = 16'b1111111110011111;
	assign R[19][13] = 16'b1111111110100100;
	assign R[19][14] = 16'b0000000001010010;
	assign R[19][15] = 16'b1111111110000000;
	assign R[19][16] = 16'b1111111110011100;
	assign R[19][17] = 16'b0000000010000010;
	assign R[19][18] = 16'b1111111111111101;
	assign R[19][19] = 16'b0000000010001000;
	assign R[19][20] = 16'b1111111111111010;
	assign R[19][21] = 16'b0000000001111110;
	assign R[19][22] = 16'b0000000000010010;
	assign R[19][23] = 16'b0000000000110001;
	assign R[19][24] = 16'b0000000000101100;
	assign R[19][25] = 16'b0000000000000111;
	assign R[19][26] = 16'b1111111111001111;
	assign R[19][27] = 16'b0000000000111000;
	assign R[19][28] = 16'b1111111110101000;
	assign R[19][29] = 16'b0000000001001010;
	assign R[19][30] = 16'b1111111111111010;
	assign R[19][31] = 16'b0000000001100011;
	assign R[20][0]  = 16'b1111111100011100;
	assign R[20][1]  = 16'b0000000000010010;
	assign R[20][2]  = 16'b1111111111111000;
	assign R[20][3]  = 16'b0000000000011010;
	assign R[20][4]  = 16'b1111111111101101;
	assign R[20][5]  = 16'b0000000001001001;
	assign R[20][6]  = 16'b0000000000000010;
	assign R[20][7]  = 16'b1111111111010110;
	assign R[20][8]  = 16'b0000000000001100;
	assign R[20][9]  = 16'b1111111110110101;
	assign R[20][10] = 16'b0000000001010101;
	assign R[20][11] = 16'b0000000000111110;
	assign R[20][12] = 16'b0000000010011111;
	assign R[20][13] = 16'b0000000001011000;
	assign R[20][14] = 16'b0000000000100000;
	assign R[20][15] = 16'b0000000000010001;
	assign R[20][16] = 16'b0000000000011101;
	assign R[20][17] = 16'b0000000000101011;
	assign R[20][18] = 16'b1111111111000000;
	assign R[20][19] = 16'b1111111110010001;
	assign R[20][20] = 16'b0000000000011001;
	assign R[20][21] = 16'b1111111111100110;
	assign R[20][22] = 16'b1111111111111011;
	assign R[20][23] = 16'b0000000000110010;
	assign R[20][24] = 16'b0000000000100011;
	assign R[20][25] = 16'b0000000000100100;
	assign R[20][26] = 16'b1111111111011011;
	assign R[20][27] = 16'b0000000010110010;
	assign R[20][28] = 16'b1111111101110110;
	assign R[20][29] = 16'b1111111101011000;
	assign R[20][30] = 16'b1111111111000110;
	assign R[20][31] = 16'b1111111110100101;
	assign R[21][0]  = 16'b1111111111001011;
	assign R[21][1]  = 16'b1111111111010101;
	assign R[21][2]  = 16'b0000000001011111;
	assign R[21][3]  = 16'b1111111110110011;
	assign R[21][4]  = 16'b0000000000101011;
	assign R[21][5]  = 16'b1111111111010110;
	assign R[21][6]  = 16'b1111111111011100;
	assign R[21][7]  = 16'b0000000000110110;
	assign R[21][8]  = 16'b0000000001001110;
	assign R[21][9]  = 16'b0000000001100110;
	assign R[21][10] = 16'b0000000000101110;
	assign R[21][11] = 16'b1111111111001001;
	assign R[21][12] = 16'b1111111111111100;
	assign R[21][13] = 16'b1111111111010011;
	assign R[21][14] = 16'b0000000000000100;
	assign R[21][15] = 16'b1111111100001011;
	assign R[21][16] = 16'b1111111110001110;
	assign R[21][17] = 16'b1111111111111111;
	assign R[21][18] = 16'b0000000000100101;
	assign R[21][19] = 16'b1111111111011001;
	assign R[21][20] = 16'b0000000000111000;
	assign R[21][21] = 16'b0000000000001000;
	assign R[21][22] = 16'b1111111111010010;
	assign R[21][23] = 16'b0000000000110101;
	assign R[21][24] = 16'b0000000000101100;
	assign R[21][25] = 16'b1111111110001110;
	assign R[21][26] = 16'b1111111110010011;
	assign R[21][27] = 16'b0000000001010010;
	assign R[21][28] = 16'b0000000010100000;
	assign R[21][29] = 16'b1111111101111000;
	assign R[21][30] = 16'b0000000000110000;
	assign R[21][31] = 16'b1111111111000001;
	assign R[22][0]  = 16'b0000000000001010;
	assign R[22][1]  = 16'b1111111111111010;
	assign R[22][2]  = 16'b0000000000011011;
	assign R[22][3]  = 16'b1111111111101100;
	assign R[22][4]  = 16'b1111111110111101;
	assign R[22][5]  = 16'b1111111111101001;
	assign R[22][6]  = 16'b1111111111011110;
	assign R[22][7]  = 16'b1111111101001000;
	assign R[22][8]  = 16'b1111111111011000;
	assign R[22][9]  = 16'b0000000000100010;
	assign R[22][10] = 16'b0000000000001000;
	assign R[22][11] = 16'b1111111111111001;
	assign R[22][12] = 16'b1111111111100111;
	assign R[22][13] = 16'b1111111110110110;
	assign R[22][14] = 16'b1111111111101011;
	assign R[22][15] = 16'b1111111110011010;
	assign R[22][16] = 16'b0000000001011001;
	assign R[22][17] = 16'b1111111111010001;
	assign R[22][18] = 16'b0000000000001111;
	assign R[22][19] = 16'b1111111111100100;
	assign R[22][20] = 16'b0000000000000010;
	assign R[22][21] = 16'b1111111111101011;
	assign R[22][22] = 16'b1111111110110000;
	assign R[22][23] = 16'b0000000000100000;
	assign R[22][24] = 16'b1111111101110101;
	assign R[22][25] = 16'b1111111110101010;
	assign R[22][26] = 16'b1111111111001100;
	assign R[22][27] = 16'b0000000000000000;
	assign R[22][28] = 16'b0000000000110001;
	assign R[22][29] = 16'b0000000000111110;
	assign R[22][30] = 16'b1111111111001111;
	assign R[22][31] = 16'b0000000000111111;
	assign R[23][0]  = 16'b0000000000111011;
	assign R[23][1]  = 16'b1111111111001001;
	assign R[23][2]  = 16'b1111111111010011;
	assign R[23][3]  = 16'b1111111111110101;
	assign R[23][4]  = 16'b0000000010110111;
	assign R[23][5]  = 16'b1111111111001001;
	assign R[23][6]  = 16'b0000000001000010;
	assign R[23][7]  = 16'b1111111111100100;
	assign R[23][8]  = 16'b0000000001000010;
	assign R[23][9]  = 16'b1111111101110101;
	assign R[23][10] = 16'b0000000001100101;
	assign R[23][11] = 16'b1111111111000011;
	assign R[23][12] = 16'b1111111111110001;
	assign R[23][13] = 16'b0000000000100010;
	assign R[23][14] = 16'b0000000000011000;
	assign R[23][15] = 16'b1111111101011010;
	assign R[23][16] = 16'b0000000000001111;
	assign R[23][17] = 16'b1111111111110100;
	assign R[23][18] = 16'b0000000000100101;
	assign R[23][19] = 16'b1111111111010111;
	assign R[23][20] = 16'b0000000001111000;
	assign R[23][21] = 16'b0000000000100010;
	assign R[23][22] = 16'b0000000010110001;
	assign R[23][23] = 16'b0000000001001101;
	assign R[23][24] = 16'b0000000000011100;
	assign R[23][25] = 16'b1111111111100111;
	assign R[23][26] = 16'b1111111101011011;
	assign R[23][27] = 16'b1111111011011111;
	assign R[23][28] = 16'b1111111111000111;
	assign R[23][29] = 16'b0000000000101001;
	assign R[23][30] = 16'b1111111111000010;
	assign R[23][31] = 16'b1111111100101110;
	assign R[24][0]  = 16'b1111111111101111;
	assign R[24][1]  = 16'b0000000001001001;
	assign R[24][2]  = 16'b0000000000000100;
	assign R[24][3]  = 16'b0000000000111110;
	assign R[24][4]  = 16'b1111111111000100;
	assign R[24][5]  = 16'b1111111110100110;
	assign R[24][6]  = 16'b0000000001000011;
	assign R[24][7]  = 16'b0000000000111000;
	assign R[24][8]  = 16'b1111111111110000;
	assign R[24][9]  = 16'b1111111111000001;
	assign R[24][10] = 16'b0000000000000001;
	assign R[24][11] = 16'b0000000000100110;
	assign R[24][12] = 16'b1111111110111100;
	assign R[24][13] = 16'b0000000001000101;
	assign R[24][14] = 16'b1111111110110001;
	assign R[24][15] = 16'b1111111111101000;
	assign R[24][16] = 16'b0000000000011110;
	assign R[24][17] = 16'b0000000000100010;
	assign R[24][18] = 16'b0000000000101100;
	assign R[24][19] = 16'b1111111111000001;
	assign R[24][20] = 16'b1111111111010111;
	assign R[24][21] = 16'b1111111111101000;
	assign R[24][22] = 16'b1111111110111110;
	assign R[24][23] = 16'b0000000000000110;
	assign R[24][24] = 16'b1111111111011001;
	assign R[24][25] = 16'b1111111111000010;
	assign R[24][26] = 16'b0000000000100000;
	assign R[24][27] = 16'b0000000001100110;
	assign R[24][28] = 16'b1111111110110010;
	assign R[24][29] = 16'b1111111110110001;
	assign R[24][30] = 16'b1111111110111110;
	assign R[24][31] = 16'b1111111110001110;
	assign R[25][0]  = 16'b0000000000011001;
	assign R[25][1]  = 16'b1111111111001001;
	assign R[25][2]  = 16'b1111111111111100;
	assign R[25][3]  = 16'b1111111110011100;
	assign R[25][4]  = 16'b1111111111001110;
	assign R[25][5]  = 16'b1111111111111000;
	assign R[25][6]  = 16'b1111111101100000;
	assign R[25][7]  = 16'b1111111101110000;
	assign R[25][8]  = 16'b1111111111100001;
	assign R[25][9]  = 16'b0000000000000000;
	assign R[25][10] = 16'b1111111111010001;
	assign R[25][11] = 16'b1111111111100000;
	assign R[25][12] = 16'b0000000010000010;
	assign R[25][13] = 16'b1111111110100011;
	assign R[25][14] = 16'b0000000000101001;
	assign R[25][15] = 16'b0000000010001101;
	assign R[25][16] = 16'b1111111111001000;
	assign R[25][17] = 16'b0000000001010101;
	assign R[25][18] = 16'b0000000000000111;
	assign R[25][19] = 16'b0000000000111101;
	assign R[25][20] = 16'b1111111111010000;
	assign R[25][21] = 16'b1111111111010001;
	assign R[25][22] = 16'b1111111100110100;
	assign R[25][23] = 16'b0000000000100100;
	assign R[25][24] = 16'b0000000001010011;
	assign R[25][25] = 16'b0000000010111011;
	assign R[25][26] = 16'b0000000000101010;
	assign R[25][27] = 16'b1111111111111010;
	assign R[25][28] = 16'b0000000001010111;
	assign R[25][29] = 16'b0000000000100010;
	assign R[25][30] = 16'b1111111110111000;
	assign R[25][31] = 16'b1111111110111101;
	assign R[26][0]  = 16'b1111111111001001;
	assign R[26][1]  = 16'b0000000000100000;
	assign R[26][2]  = 16'b0000000000111111;
	assign R[26][3]  = 16'b1111111111110100;
	assign R[26][4]  = 16'b1111111110100010;
	assign R[26][5]  = 16'b0000000000000010;
	assign R[26][6]  = 16'b1111111111011111;
	assign R[26][7]  = 16'b1111111110000011;
	assign R[26][8]  = 16'b0000000000001010;
	assign R[26][9]  = 16'b1111111111101001;
	assign R[26][10] = 16'b0000000001111110;
	assign R[26][11] = 16'b1111111111100110;
	assign R[26][12] = 16'b0000000000010100;
	assign R[26][13] = 16'b0000000000111010;
	assign R[26][14] = 16'b0000000000010000;
	assign R[26][15] = 16'b1111111111001011;
	assign R[26][16] = 16'b0000000000001000;
	assign R[26][17] = 16'b1111111111011111;
	assign R[26][18] = 16'b1111111110011000;
	assign R[26][19] = 16'b1111111110111101;
	assign R[26][20] = 16'b0000000000101011;
	assign R[26][21] = 16'b0000000001001100;
	assign R[26][22] = 16'b1111111110101100;
	assign R[26][23] = 16'b0000000010000001;
	assign R[26][24] = 16'b0000000000010111;
	assign R[26][25] = 16'b1111111110001001;
	assign R[26][26] = 16'b1111111110111111;
	assign R[26][27] = 16'b1111111111101111;
	assign R[26][28] = 16'b0000000000111010;
	assign R[26][29] = 16'b1111111110000001;
	assign R[26][30] = 16'b1111111111010110;
	assign R[26][31] = 16'b0000000000110100;
	assign R[27][0]  = 16'b0000000000001010;
	assign R[27][1]  = 16'b0000000010000000;
	assign R[27][2]  = 16'b0000000000011101;
	assign R[27][3]  = 16'b0000000000011110;
	assign R[27][4]  = 16'b1111111111010110;
	assign R[27][5]  = 16'b0000000000010110;
	assign R[27][6]  = 16'b0000000010001000;
	assign R[27][7]  = 16'b1111111111111011;
	assign R[27][8]  = 16'b1111111111010010;
	assign R[27][9]  = 16'b0000000000101100;
	assign R[27][10] = 16'b1111111111100110;
	assign R[27][11] = 16'b0000000000111010;
	assign R[27][12] = 16'b0000000010100001;
	assign R[27][13] = 16'b1111111111001000;
	assign R[27][14] = 16'b0000000000111000;
	assign R[27][15] = 16'b0000000001111101;
	assign R[27][16] = 16'b0000000000001111;
	assign R[27][17] = 16'b0000000000001111;
	assign R[27][18] = 16'b0000000010010011;
	assign R[27][19] = 16'b1111111111110011;
	assign R[27][20] = 16'b1111111111010101;
	assign R[27][21] = 16'b1111111111011011;
	assign R[27][22] = 16'b1111111110011011;
	assign R[27][23] = 16'b1111111111100110;
	assign R[27][24] = 16'b1111111111011110;
	assign R[27][25] = 16'b0000000000111101;
	assign R[27][26] = 16'b0000000001000110;
	assign R[27][27] = 16'b1111111110111011;
	assign R[27][28] = 16'b1111111111100100;
	assign R[27][29] = 16'b1111111110111100;
	assign R[27][30] = 16'b0000000000011100;
	assign R[27][31] = 16'b1111111111110000;
	assign R[28][0]  = 16'b0000000000011111;
	assign R[28][1]  = 16'b1111111110011000;
	assign R[28][2]  = 16'b1111111111101000;
	assign R[28][3]  = 16'b1111111111100110;
	assign R[28][4]  = 16'b1111111111010001;
	assign R[28][5]  = 16'b1111111111000110;
	assign R[28][6]  = 16'b1111111111001001;
	assign R[28][7]  = 16'b0000000000011100;
	assign R[28][8]  = 16'b0000000000101111;
	assign R[28][9]  = 16'b0000000001001000;
	assign R[28][10] = 16'b1111111111110101;
	assign R[28][11] = 16'b1111111110110100;
	assign R[28][12] = 16'b0000000000011001;
	assign R[28][13] = 16'b1111111110011000;
	assign R[28][14] = 16'b1111111110111011;
	assign R[28][15] = 16'b1111111101000100;
	assign R[28][16] = 16'b1111111101100110;
	assign R[28][17] = 16'b1111111110010111;
	assign R[28][18] = 16'b1111111110100100;
	assign R[28][19] = 16'b1111111111010010;
	assign R[28][20] = 16'b1111111111110101;
	assign R[28][21] = 16'b0000000000101011;
	assign R[28][22] = 16'b1111111110111000;
	assign R[28][23] = 16'b1111111111011111;
	assign R[28][24] = 16'b1111111101110011;
	assign R[28][25] = 16'b0000000000011001;
	assign R[28][26] = 16'b0000000000101011;
	assign R[28][27] = 16'b0000000001100001;
	assign R[28][28] = 16'b0000000000100001;
	assign R[28][29] = 16'b1111111111000100;
	assign R[28][30] = 16'b1111111111101010;
	assign R[28][31] = 16'b0000000000001011;
	assign R[29][0]  = 16'b1111111110011111;
	assign R[29][1]  = 16'b0000000001001000;
	assign R[29][2]  = 16'b0000000000100000;
	assign R[29][3]  = 16'b0000000001101101;
	assign R[29][4]  = 16'b1111111111011101;
	assign R[29][5]  = 16'b0000000001100010;
	assign R[29][6]  = 16'b1111111101111110;
	assign R[29][7]  = 16'b0000000001101000;
	assign R[29][8]  = 16'b0000000001001101;
	assign R[29][9]  = 16'b0000000001110011;
	assign R[29][10] = 16'b0000000000100101;
	assign R[29][11] = 16'b0000000000011101;
	assign R[29][12] = 16'b1111111111111010;
	assign R[29][13] = 16'b0000000001110011;
	assign R[29][14] = 16'b0000000000010110;
	assign R[29][15] = 16'b0000000000101101;
	assign R[29][16] = 16'b0000000000101001;
	assign R[29][17] = 16'b1111111111111100;
	assign R[29][18] = 16'b1111111110101100;
	assign R[29][19] = 16'b0000000000000110;
	assign R[29][20] = 16'b0000000000111111;
	assign R[29][21] = 16'b1111111110111110;
	assign R[29][22] = 16'b0000000000010110;
	assign R[29][23] = 16'b0000000001100111;
	assign R[29][24] = 16'b0000000000001100;
	assign R[29][25] = 16'b1111111111011100;
	assign R[29][26] = 16'b0000000000110111;
	assign R[29][27] = 16'b0000000001101101;
	assign R[29][28] = 16'b0000000001001001;
	assign R[29][29] = 16'b0000000000110100;
	assign R[29][30] = 16'b1111111111001001;
	assign R[29][31] = 16'b0000000010001001;
	assign R[30][0]  = 16'b1111111111010110;
	assign R[30][1]  = 16'b0000000000011111;
	assign R[30][2]  = 16'b0000000000000011;
	assign R[30][3]  = 16'b0000000000000000;
	assign R[30][4]  = 16'b1111111111111001;
	assign R[30][5]  = 16'b1111111111100000;
	assign R[30][6]  = 16'b0000000000001000;
	assign R[30][7]  = 16'b1111111111011100;
	assign R[30][8]  = 16'b1111111111110000;
	assign R[30][9]  = 16'b1111111111110000;
	assign R[30][10] = 16'b1111111111101011;
	assign R[30][11] = 16'b1111111111000001;
	assign R[30][12] = 16'b0000000001111110;
	assign R[30][13] = 16'b0000000000001001;
	assign R[30][14] = 16'b0000000001001011;
	assign R[30][15] = 16'b1111111111110111;
	assign R[30][16] = 16'b0000000001101111;
	assign R[30][17] = 16'b1111111111110111;
	assign R[30][18] = 16'b0000000000110111;
	assign R[30][19] = 16'b1111111101111010;
	assign R[30][20] = 16'b1111111111011000;
	assign R[30][21] = 16'b1111111111101101;
	assign R[30][22] = 16'b1111111110111000;
	assign R[30][23] = 16'b0000000000101100;
	assign R[30][24] = 16'b1111111110001101;
	assign R[30][25] = 16'b0000000001000101;
	assign R[30][26] = 16'b0000000001001101;
	assign R[30][27] = 16'b1111111111101110;
	assign R[30][28] = 16'b0000000001010011;
	assign R[30][29] = 16'b1111111110110101;
	assign R[30][30] = 16'b0000000011011111;
	assign R[30][31] = 16'b1111111100010101;
	assign R[31][0]  = 16'b0000000001011000;
	assign R[31][1]  = 16'b1111111111011011;
	assign R[31][2]  = 16'b1111111110111110;
	assign R[31][3]  = 16'b1111111110111001;
	assign R[31][4]  = 16'b0000000000011001;
	assign R[31][5]  = 16'b0000000000000010;
	assign R[31][6]  = 16'b1111111110111001;
	assign R[31][7]  = 16'b1111111111001000;
	assign R[31][8]  = 16'b0000000000110010;
	assign R[31][9]  = 16'b1111111111100001;
	assign R[31][10] = 16'b1111111110100011;
	assign R[31][11] = 16'b1111111111110000;
	assign R[31][12] = 16'b0000000000001101;
	assign R[31][13] = 16'b0000000000100010;
	assign R[31][14] = 16'b1111111111010011;
	assign R[31][15] = 16'b0000000001011111;
	assign R[31][16] = 16'b1111111110001101;
	assign R[31][17] = 16'b0000000010011001;
	assign R[31][18] = 16'b0000000001010110;
	assign R[31][19] = 16'b0000000000001011;
	assign R[31][20] = 16'b0000000000011001;
	assign R[31][21] = 16'b0000000001010110;
	assign R[31][22] = 16'b0000000000011100;
	assign R[31][23] = 16'b0000000000001000;
	assign R[31][24] = 16'b1111111111100011;
	assign R[31][25] = 16'b0000000000010011;
	assign R[31][26] = 16'b1111111111110000;
	assign R[31][27] = 16'b0000000001110111;
	assign R[31][28] = 16'b1111111101101000;
	assign R[31][29] = 16'b1111111111011010;
	assign R[31][30] = 16'b0000000000010100;
	assign R[31][31] = 16'b1111111111000111;

endmodule