module rnn_bias();

	logic [15:0] RB[0:31];

	assign RB[0 ] = 16'b1111111111000001;
	assign RB[1 ] = 16'b1111111111011000;
	assign RB[2 ] = 16'b1111111101100001;
	assign RB[3 ] = 16'b1111111111101011;
	assign RB[4 ] = 16'b0000000001100111;
	assign RB[5 ] = 16'b1111111111000000;
	assign RB[6 ] = 16'b0000000010011010;
	assign RB[7 ] = 16'b1111111010100011;
	assign RB[8 ] = 16'b0000000000001100;
	assign RB[9 ] = 16'b0000000000000000;
	assign RB[10] = 16'b0000000001000000;
	assign RB[11] = 16'b0000000000101110;
	assign RB[12] = 16'b0000000000001001;
	assign RB[13] = 16'b0000000000111110;
	assign RB[14] = 16'b0000000000110111;
	assign RB[15] = 16'b1111111111001101;
	assign RB[16] = 16'b1111111110000111;
	assign RB[17] = 16'b0000000000100110;
	assign RB[18] = 16'b0000000001110001;
	assign RB[19] = 16'b0000000000101101;
	assign RB[20] = 16'b1111111111000010;
	assign RB[21] = 16'b0000000010001111;
	assign RB[22] = 16'b0000000011110101;
	assign RB[23] = 16'b0000000001010110;
	assign RB[24] = 16'b1111111111001111;
	assign RB[25] = 16'b1111111110100110;
	assign RB[26] = 16'b1111111111010111;
	assign RB[27] = 16'b1111111110000111;
	assign RB[28] = 16'b1111111110101010;
	assign RB[29] = 16'b1111111101100010;
	assign RB[30] = 16'b0000000000100001;
	assign RB[31] = 16'b1111111111000011;

endmodule : rnn_bias