module tanh_tb();

	logic signed [15:0] in, out, guess, difference;
	tanh dut(.*);

assign difference = (guess - out) >= 0 ? guess - out: out - guess;

// automatically generated testbench using python
// tests for a range of fixed point values ranging from -2 to 2 in increments of 0.1

	initial begin
in = 16'b11111100_00000000;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_00011010;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_00110100;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_01001101;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_01100111;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_10000000;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_10011010;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_10110100;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_11001101;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111100_11100111;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_00000000;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_00011010;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_00110100;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_01001101;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_01100111;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_10000000;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_10011010;
guess = 16'b11111111_00000000;
assert(difference <= 1);
#5;
in = 16'b11111101_10110100;
guess = 16'b11111111_00000100;
assert(difference <= 1);
#5;
in = 16'b11111101_11001101;
guess = 16'b11111111_00000111;
assert(difference <= 1);
#5;
in = 16'b11111101_11100111;
guess = 16'b11111111_00001010;
assert(difference <= 1);
#5;
in = 16'b11111110_00000000;
guess = 16'b11111111_00001101;
assert(difference <= 1);
#5;
in = 16'b11111110_00011010;
guess = 16'b11111111_00010000;
assert(difference <= 1);
#5;
in = 16'b11111110_00110100;
guess = 16'b11111111_00010100;
assert(difference <= 1);
#5;
in = 16'b11111110_01001101;
guess = 16'b11111111_00010111;
assert(difference <= 1);
#5;
in = 16'b11111110_01100111;
guess = 16'b11111111_00011010;
assert(difference <= 1);
#5;
in = 16'b11111110_10000000;
guess = 16'b11111111_00011101;
assert(difference <= 1);
#5;
in = 16'b11111110_10011010;
guess = 16'b11111111_00100000;
assert(difference <= 1);
#5;
in = 16'b11111110_10110100;
guess = 16'b11111111_00100100;
assert(difference <= 1);
#5;
in = 16'b11111110_11001101;
guess = 16'b11111111_00100111;
assert(difference <= 1);
#5;
in = 16'b11111110_11100111;
guess = 16'b11111111_00110100;
assert(difference <= 1);
#5;
in = 16'b11111111_00000000;
guess = 16'b11111111_01000000;
assert(difference <= 1);
#5;
in = 16'b11111111_00011010;
guess = 16'b11111111_01001101;
assert(difference <= 1);
#5;
in = 16'b11111111_00110100;
guess = 16'b11111111_01011010;
assert(difference <= 1);
#5;
in = 16'b11111111_01001101;
guess = 16'b11111111_01100111;
assert(difference <= 1);
#5;
in = 16'b11111111_01100111;
guess = 16'b11111111_01110100;
assert(difference <= 1);
#5;
in = 16'b11111111_10000000;
guess = 16'b11111111_10000000;
assert(difference <= 1);
#5;
in = 16'b11111111_10011010;
guess = 16'b11111111_10011010;
assert(difference <= 1);
#5;
in = 16'b11111111_10110100;
guess = 16'b11111111_10110100;
assert(difference <= 1);
#5;
in = 16'b11111111_11001101;
guess = 16'b11111111_11001101;
assert(difference <= 1);
#5;
in = 16'b11111111_11100111;
guess = 16'b11111111_11100111;
assert(difference <= 1);
#5;
in = 16'b00000000_00000000;
guess = 16'b00000000_00000000;
assert(difference <= 1);
#5;
in = 16'b00000000_00011001;
guess = 16'b00000000_00011001;
assert(difference <= 1);
#5;
in = 16'b00000000_00110011;
guess = 16'b00000000_00110011;
assert(difference <= 1);
#5;
in = 16'b00000000_01001100;
guess = 16'b00000000_01001100;
assert(difference <= 1);
#5;
in = 16'b00000000_01100110;
guess = 16'b00000000_01100110;
assert(difference <= 1);
#5;
in = 16'b00000000_10000000;
guess = 16'b00000000_10000000;
assert(difference <= 1);
#5;
in = 16'b00000000_10011001;
guess = 16'b00000000_10001100;
assert(difference <= 1);
#5;
in = 16'b00000000_10110011;
guess = 16'b00000000_10011001;
assert(difference <= 1);
#5;
in = 16'b00000000_11001100;
guess = 16'b00000000_10100110;
assert(difference <= 1);
#5;
in = 16'b00000000_11100110;
guess = 16'b00000000_10110011;
assert(difference <= 1);
#5;
in = 16'b00000001_00000000;
guess = 16'b00000000_11000000;
assert(difference <= 1);
#5;
in = 16'b00000001_00011001;
guess = 16'b00000000_11001100;
assert(difference <= 1);
#5;
in = 16'b00000001_00110011;
guess = 16'b00000000_11011001;
assert(difference <= 1);
#5;
in = 16'b00000001_01001100;
guess = 16'b00000000_11011100;
assert(difference <= 1);
#5;
in = 16'b00000001_01100110;
guess = 16'b00000000_11100000;
assert(difference <= 1);
#5;
in = 16'b00000001_10000000;
guess = 16'b00000000_11100011;
assert(difference <= 1);
#5;
in = 16'b00000001_10011001;
guess = 16'b00000000_11100110;
assert(difference <= 1);
#5;
in = 16'b00000001_10110011;
guess = 16'b00000000_11101001;
assert(difference <= 1);
#5;
in = 16'b00000001_11001100;
guess = 16'b00000000_11101100;
assert(difference <= 1);
#5;
in = 16'b00000001_11100110;
guess = 16'b00000000_11110000;
assert(difference <= 1);
#5;
in = 16'b00000010_00000000;
guess = 16'b00000000_11110011;
assert(difference <= 1);
#5;
in = 16'b00000010_00011001;
guess = 16'b00000000_11110110;
assert(difference <= 1);
#5;
in = 16'b00000010_00110011;
guess = 16'b00000000_11111001;
assert(difference <= 1);
#5;
in = 16'b00000010_01001100;
guess = 16'b00000000_11111100;
assert(difference <= 1);
#5;
in = 16'b00000010_01100110;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000010_10000000;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000010_10011001;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000010_10110011;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000010_11001100;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000010_11100110;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_00000000;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_00011001;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_00110011;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_01001100;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_01100110;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_10000000;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_10011001;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_10110011;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_11001100;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;
in = 16'b00000011_11100110;
guess = 16'b00000001_00000000;
assert(difference <= 1);
#5;

	end
endmodule