module dense();

	logic [15:0] D[0:31];

	assign D[0 ] = 16'b0000000000111100;
	assign D[1 ] = 16'b1111111110100000;
	assign D[2 ] = 16'b1111111110001000;
	assign D[3 ] = 16'b1111111101111011;
	assign D[4 ] = 16'b0000000011000100;
	assign D[5 ] = 16'b0000000001101101;
	assign D[6 ] = 16'b0000000000011101;
	assign D[7 ] = 16'b0000000000011110;
	assign D[8 ] = 16'b0000000010100100;
	assign D[9 ] = 16'b1111111111111110;
	assign D[10] = 16'b0000000000000110;
	assign D[11] = 16'b1111111110010010;
	assign D[12] = 16'b1111111111100101;
	assign D[13] = 16'b0000000010111111;
	assign D[14] = 16'b1111111111110010;
	assign D[15] = 16'b0000000000001111;
	assign D[16] = 16'b1111111101111111;
	assign D[17] = 16'b0000000000010000;
	assign D[18] = 16'b1111111110100001;
	assign D[19] = 16'b0000000000101010;
	assign D[20] = 16'b0000000010110101;
	assign D[21] = 16'b0000000010001010;
	assign D[22] = 16'b0000000001100101;
	assign D[23] = 16'b0000000000110110;
	assign D[24] = 16'b1111111111001100;
	assign D[25] = 16'b1111111111001010;
	assign D[26] = 16'b1111111101001011;
	assign D[27] = 16'b0000000000001011;
	assign D[28] = 16'b1111111110000001;
	assign D[29] = 16'b0000000001011110;
	assign D[30] = 16'b1111111110001001;
	assign D[31] = 16'b0000000000101111;

endmodule