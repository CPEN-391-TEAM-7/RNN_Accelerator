
module rnn(
	input  logic clk,
	input  logic rst_n
	);



endmodule : rnn