module embedding();

	logic [15:0] E[0:38][0:3];
	
	assign E[0][0]  = 16'b1111111110001111;
 	assign E[0][1]  = 16'b0000000110110011;
 	assign E[0][2]  = 16'b1111111101000001;
 	assign E[0][3]  = 16'b0000000001001111;
 	assign E[1][0]  = 16'b1111111100001000;
 	assign E[1][1]  = 16'b1111111101110000;
 	assign E[1][2]  = 16'b0000000001101000;
 	assign E[1][3]  = 16'b0000000000000101;
 	assign E[2][0]  = 16'b0000000010010111;
 	assign E[2][1]  = 16'b1111111110001010;
 	assign E[2][2]  = 16'b1111111110111111;
 	assign E[2][3]  = 16'b1111111110101110;
 	assign E[3][0]  = 16'b1111111011100001;
 	assign E[3][1]  = 16'b1111111111100010;
 	assign E[3][2]  = 16'b0000000001001000;
 	assign E[3][3]  = 16'b0000000000000000;
 	assign E[4][0]  = 16'b1111111111101100;
 	assign E[4][1]  = 16'b0000000001001001;
 	assign E[4][2]  = 16'b1111111110000110;
 	assign E[4][3]  = 16'b0000000001011101;
 	assign E[5][0]  = 16'b1111111010110000;
 	assign E[5][1]  = 16'b1111111101000010;
 	assign E[5][2]  = 16'b0000000000111111;
 	assign E[5][3]  = 16'b0000000000111001;
 	assign E[6][0]  = 16'b1111111011110100;
 	assign E[6][1]  = 16'b1111111110010101;
 	assign E[6][2]  = 16'b0000000000101011;
 	assign E[6][3]  = 16'b0000000000001100;
 	assign E[7][0]  = 16'b1111111111000101;
 	assign E[7][1]  = 16'b1111111110011011;
 	assign E[7][2]  = 16'b0000000000011011;
 	assign E[7][3]  = 16'b0000000000000000;
 	assign E[8][0]  = 16'b0000000001001001;
 	assign E[8][1]  = 16'b0000000000110011;
 	assign E[8][2]  = 16'b1111111110100100;
 	assign E[8][3]  = 16'b0000000001101100;
 	assign E[9][0]  = 16'b1111111101000000;
 	assign E[9][1]  = 16'b1111111001111001;
 	assign E[9][2]  = 16'b0000000000111100;
 	assign E[9][3]  = 16'b1111111111100110;
 	assign E[10][0] = 16'b1111111001100010;
 	assign E[10][1] = 16'b1111111101110000;
 	assign E[10][2] = 16'b0000000001010010;
 	assign E[10][3] = 16'b0000000001000101;
 	assign E[11][0] = 16'b1111111011010011;
 	assign E[11][1] = 16'b0000000000001101;
 	assign E[11][2] = 16'b0000000010101000;
 	assign E[11][3] = 16'b0000000000111000;
 	assign E[12][0] = 16'b1111111101101111;
 	assign E[12][1] = 16'b1111111110011100;
 	assign E[12][2] = 16'b1111111111110111;
 	assign E[12][3] = 16'b1111111111011000;
 	assign E[13][0] = 16'b1111111100001101;
 	assign E[13][1] = 16'b1111111110101010;
 	assign E[13][2] = 16'b0000000011100101;
 	assign E[13][3] = 16'b0000000001111111;
 	assign E[14][0] = 16'b1111111111101010;
 	assign E[14][1] = 16'b0000000001101111;
 	assign E[14][2] = 16'b1111111110000010;
 	assign E[14][3] = 16'b0000000001011001;
 	assign E[15][0] = 16'b1111111001011100;
 	assign E[15][1] = 16'b1111111111010111;
 	assign E[15][2] = 16'b0000000000111001;
 	assign E[15][3] = 16'b0000000001001001;
 	assign E[16][0] = 16'b1111110101110100;
 	assign E[16][1] = 16'b1111110111100000;
 	assign E[16][2] = 16'b0000000001011001;
 	assign E[16][3] = 16'b0000000000100100;
 	assign E[17][0] = 16'b1111111100100110;
 	assign E[17][1] = 16'b0000000000110010;
 	assign E[17][2] = 16'b0000000010010001;
 	assign E[17][3] = 16'b0000000000111001;
 	assign E[18][0] = 16'b1111111011111100;
 	assign E[18][1] = 16'b0000000010110101;
 	assign E[18][2] = 16'b1111111111011001;
 	assign E[18][3] = 16'b0000000000000011;
 	assign E[19][0] = 16'b1111111010010101;
 	assign E[19][1] = 16'b0000000001011110;
 	assign E[19][2] = 16'b0000000001010100;
 	assign E[19][3] = 16'b0000000000101010;
 	assign E[20][0] = 16'b0000000001000111;
 	assign E[20][1] = 16'b1111111110011011;
 	assign E[20][2] = 16'b1111111101100110;
 	assign E[20][3] = 16'b0000000000101100;
 	assign E[21][0] = 16'b1111111001011101;
 	assign E[21][1] = 16'b1111111100100010;
 	assign E[21][2] = 16'b0000000001101001;
 	assign E[21][3] = 16'b0000000000100110;
 	assign E[22][0] = 16'b1111111111100001;
 	assign E[22][1] = 16'b1111111010101100;
 	assign E[22][2] = 16'b0000000000000011;
 	assign E[22][3] = 16'b1111111111101010;
 	assign E[23][0] = 16'b1111111101000110;
 	assign E[23][1] = 16'b1111111010101100;
 	assign E[23][2] = 16'b0000000000001110;
 	assign E[23][3] = 16'b1111111111011110;
 	assign E[24][0] = 16'b1111111100000110;
 	assign E[24][1] = 16'b0000000000001100;
 	assign E[24][2] = 16'b1111111100100000;
 	assign E[24][3] = 16'b1111111111101000;
 	assign E[25][0] = 16'b1111111101110001;
 	assign E[25][1] = 16'b1111111110001000;
 	assign E[25][2] = 16'b0000000000011011;
 	assign E[25][3] = 16'b0000000000000011;
 	assign E[26][0] = 16'b1111111100101011;
 	assign E[26][1] = 16'b0000001011110111;
 	assign E[26][2] = 16'b1111111101110110;
 	assign E[26][3] = 16'b1111111111011010;
 	assign E[27][0] = 16'b0000000000101110;
 	assign E[27][1] = 16'b1111111100110011;
 	assign E[27][2] = 16'b1111111101001011;
 	assign E[27][3] = 16'b1111111100000000;
 	assign E[28][0] = 16'b0000000000101101;
 	assign E[28][1] = 16'b1111111111010110;
 	assign E[28][2] = 16'b1111111100101101;
 	assign E[28][3] = 16'b1111111101000001;
 	assign E[29][0] = 16'b0000000000010101;
 	assign E[29][1] = 16'b1111111011010101;
 	assign E[29][2] = 16'b1111111101011011;
 	assign E[29][3] = 16'b1111111100001110;
 	assign E[30][0] = 16'b0000000001001101;
 	assign E[30][1] = 16'b1111111100111101;
 	assign E[30][2] = 16'b1111111100101111;
 	assign E[30][3] = 16'b1111111100010001;
 	assign E[31][0] = 16'b0000000000000000;
 	assign E[31][1] = 16'b1111111000111111;
 	assign E[31][2] = 16'b1111111101101100;
 	assign E[31][3] = 16'b1111111011110010;
 	assign E[32][0] = 16'b1111111111111100;
 	assign E[32][1] = 16'b1111110111111101;
 	assign E[32][2] = 16'b1111111101101000;
 	assign E[32][3] = 16'b1111111011101001;
 	assign E[33][0] = 16'b1111111111110111;
 	assign E[33][1] = 16'b1111111001100011;
 	assign E[33][2] = 16'b1111111101101001;
 	assign E[33][3] = 16'b1111111100000110;
 	assign E[34][0] = 16'b1111111111101001;
 	assign E[34][1] = 16'b1111111000110010;
 	assign E[34][2] = 16'b1111111101100011;
 	assign E[34][3] = 16'b1111111010111111;
 	assign E[35][0] = 16'b1111111111100011;
 	assign E[35][1] = 16'b1111111011001100;
 	assign E[35][2] = 16'b1111111101111110;
 	assign E[35][3] = 16'b1111111011101010;
 	assign E[36][0] = 16'b0000000111101011;
 	assign E[36][1] = 16'b0000000111101001;
 	assign E[36][2] = 16'b0000000110110011;
 	assign E[36][3] = 16'b0000000100011101;
 	assign E[37][0] = 16'b1111111111111010;
 	assign E[37][1] = 16'b0000100101011001;
 	assign E[37][2] = 16'b1111111100000110;
 	assign E[37][3] = 16'b0000000001001000;
 	assign E[38][0] = 16'b1111111111111110;
 	assign E[38][1] = 16'b1111111111110111;
 	assign E[38][2] = 16'b0000000000001000;
 	assign E[38][3] = 16'b0000000000001100;

 endmodule